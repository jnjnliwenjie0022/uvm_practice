`ifndef MY_ENV__SV
`define MY_ENV__SV

class my_env extends uvm_env;
    my_agent  i_agt;
    my_agent  o_agt;
    my_model  mdl;
    uvm_tlm_analysis_fifo #(my_transaction) agt_mdl_fifo;
    my_scoreboard scb;
    uvm_tlm_analysis_fifo #(my_transaction) agt_scb_fifo;
    uvm_tlm_analysis_fifo #(my_transaction) mdl_scb_fifo;
    `uvm_component_utils(my_env)
    function new(string name = "my_env", uvm_component parent);
        super.new(name, parent);
    endfunction

    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        i_agt = my_agent::type_id::create("i_agt", this);
        o_agt = my_agent::type_id::create("o_agt", this);
        i_agt.is_active = UVM_ACTIVE;
        o_agt.is_active = UVM_PASSIVE; 
        mdl = my_model::type_id::create("mdl", this);
        agt_mdl_fifo = new("agt_mdl_fifo", this);
        scb = my_scoreboard::type_id::create("scb", this);
        agt_scb_fifo = new("agt_scb_fifo", this);
        mdl_scb_fifo = new("mdl_scb_fifo", this);
        //uvm_config_db#(uvm_object_wrapper)::set(this,
        //                                       "i_agt.sqr.main_phase",
        //                                       "default_sequence",
        //                                        my_sequence::type_id::get());
    endfunction


    extern virtual function void connect_phase(uvm_phase phase);
    //extern virtual task main_phase(uvm_phase phase);
endclass

function void my_env::connect_phase(uvm_phase phase);
    super.connect_phase(phase);
    i_agt.ap.connect(agt_mdl_fifo.analysis_export);
    mdl.port.connect(agt_mdl_fifo.blocking_get_export);
    mdl.ap.connect(mdl_scb_fifo.analysis_export);
    scb.exp_port.connect(mdl_scb_fifo.blocking_get_export);
    o_agt.ap.connect(agt_scb_fifo.analysis_export);
    scb.act_port.connect(agt_scb_fifo.blocking_get_export); 
endfunction
//task my_env::main_phase(uvm_phase phase);
//   my_sequence seq;
//   phase.raise_objection(this);
//   seq = my_sequence::type_id::create("seq");
//   seq.start(i_agt.sqr); 
//   phase.drop_objection(this);
//endtask
`endif
