`ifndef MY_MONITOR__SV
`define MY_MONITOR__SV
class my_monitor extends uvm_monitor;

    virtual my_if vif;
    //{{{
    uvm_analysis_port #(my_transaction)  ap;
    //}}}
    `uvm_component_utils(my_monitor)
    function new(string name = "my_monitor", uvm_component parent = null);
        super.new(name, parent);
    endfunction

    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        if(!uvm_config_db#(virtual my_if)::get(this, "", "vif", vif))
            `uvm_fatal("my_monitor", "virtual interface must be set for vif!!!")
        //{{{
        ap = new("ap", this);
        //}}}
    endfunction

    extern task run_phase(uvm_phase phase);
    extern task collect_one_pkt(my_transaction tr);
endclass

task my_monitor::run_phase(uvm_phase phase);
    my_transaction tr;
    while(1) begin
        tr = new("tr");
        collect_one_pkt(tr);
        `uvm_info(get_type_name(), $sformatf("Contents: \n%s", tr.sprint()), UVM_LOW)
        //{{{
        ap.write(tr);
        //}}}
    end
endtask

task my_monitor::collect_one_pkt(my_transaction tr);
   //bit[7:0] data_q[$];
   //int psize;

   byte unsigned data_q[$];
   byte unsigned data_array[];
   logic [7:0] data;
   logic valid = 0;
   int data_size;

   while(1) begin
      @(posedge vif.clk);
      if(vif.valid) break;
   end

   `uvm_info("my_monitor", "begin to collect one pkt", UVM_LOW);
   while(vif.valid) begin
      data_q.push_back(vif.data);
      @(posedge vif.clk);
   end
   ////pop dmac
   //for(int i = 0; i < 6; i++) begin
   //   tr.dmac = {tr.dmac[39:0], data_q.pop_front()};
   //end
   ////pop smac
   //for(int i = 0; i < 6; i++) begin
   //   tr.smac = {tr.smac[39:0], data_q.pop_front()};
   //end
   ////pop ether_type
   //for(int i = 0; i < 2; i++) begin
   //   tr.ether_type = {tr.ether_type[7:0], data_q.pop_front()};
   //end

   //psize = data_q.size() - 4;
   //tr.pload = new[psize];
   ////pop payload
   //for(int i = 0; i < psize; i++) begin
   //   tr.pload[i] = data_q.pop_front();
   //end
   ////pop crc
   //for(int i = 0; i < 4; i++) begin
   //   tr.crc = {tr.crc[23:0], data_q.pop_front()};
   //end
   //`uvm_info("my_monitor", "end collect one pkt, print it:", UVM_LOW);
   //tr.my_print();
   data_size  = data_q.size();
   data_array = new[data_size];
   for ( int i = 0; i < data_size; i++ ) begin
      data_array[i] = data_q[i];
   end
   tr.pload = new[data_size - 20]; //da, sa, e_type, crc
   data_size = tr.unpack_bytes(data_array) / 8;
   //data_size = tr.unpack_bytes(data_q) / 8;
   `uvm_info("my_monitor", "end collect one pkt", UVM_LOW);

endtask


`endif
